// Camera_Interface.v

// Generated using ACDS version 13.0sp1 232 at 2015.02.18.18:49:44

`timescale 1 ps / 1 ps
module Camera_Interface (
		input  wire  clk_clk,       //   clk.clk
		input  wire  reset_reset_n  // reset.reset_n
	);

	CCD_avalon_interface trdb_d5m_camera_0 (
		.iclk        (clk_clk), //   iCLK_sink.clk
		.odval       (),        //       odval.export
		.iswitches   (),        //   iswitches.export
		.ikeys       (),        //       ikeys.export
		.ored        (),        //        orgb.export
		.ogreen      (),        //            .export
		.oblue       (),        //            .export
		.oy_cont     (),        //     oy_cont.export
		.omem_rst    (),        //    omem_rst.reset
		.ovga_rst    (),        //    ovga_rst.reset
		.iogpio      (),        //      iogpio.export
		.oframe_cont (),        // oframe_cont.export
		.opixclk     (),        //     opixclk.clk
		.orclk       ()         //       orclk.export
	);

endmodule
