// Camera_Interface.v

// Generated using ACDS version 13.0sp1 232 at 2015.02.17.16:54:55

`timescale 1 ps / 1 ps
module Camera_Interface (
		input  wire        clk_clk,                                  //                                 clk.clk
		input  wire        reset_reset_n,                            //                               reset.reset_n
		input  wire        trdb_d5m_camera_0_ccd_pixclk_clk,         //        trdb_d5m_camera_0_ccd_pixclk.clk
		output wire        trdb_d5m_camera_0_orst_0_reset,           //            trdb_d5m_camera_0_orst_0.reset
		output wire        trdb_d5m_camera_0_orst_2_reset,           //            trdb_d5m_camera_0_orst_2.reset
		output wire        trdb_d5m_camera_0_orst_1_reset,           //            trdb_d5m_camera_0_orst_1.reset
		input  wire [11:0] trdb_d5m_camera_0_idata_export,           //             trdb_d5m_camera_0_idata.export
		input  wire        trdb_d5m_camera_0_iend_export,            //              trdb_d5m_camera_0_iend.export
		input  wire        trdb_d5m_camera_0_iflval_ifval,           //            trdb_d5m_camera_0_iflval.ifval
		input  wire        trdb_d5m_camera_0_iflval_ilval,           //                                    .ilval
		input  wire        trdb_d5m_camera_0_istart_export,          //            trdb_d5m_camera_0_istart.export
		input  wire        trdb_d5m_camera_0_zoom_mode_export,       //         trdb_d5m_camera_0_zoom_mode.export
		output wire [11:0] trdb_d5m_camera_0_rgb_ored,               //               trdb_d5m_camera_0_rgb.ored
		output wire [11:0] trdb_d5m_camera_0_rgb_ogreen,             //                                    .ogreen
		output wire [11:0] trdb_d5m_camera_0_rgb_oblue,              //                                    .oblue
		output wire        trdb_d5m_camera_0_odval_export,           //             trdb_d5m_camera_0_odval.export
		output wire [15:0] trdb_d5m_camera_0_oycont_export,          //            trdb_d5m_camera_0_oycont.export
		output wire [31:0] trdb_d5m_camera_0_oframe_export,          //            trdb_d5m_camera_0_oframe.export
		input  wire        trdb_d5m_camera_0_exposure_adjust_adj,    //   trdb_d5m_camera_0_exposure_adjust.adj
		input  wire        trdb_d5m_camera_0_exposure_adjust_dec_p,  //                                    .dec_p
		output wire        trdb_d5m_camera_0_i2c_configuration_sclk, // trdb_d5m_camera_0_i2c_configuration.sclk
		output wire        trdb_d5m_camera_0_i2c_configuration_sdat  //                                    .sdat
	);

	wire    rst_controller_reset_out_reset; // rst_controller:reset_out -> TRDB_D5M_Camera_0:irst

	CCD_avalon_interface trdb_d5m_camera_0 (
		.i2c_sclk        (trdb_d5m_camera_0_i2c_configuration_sclk), // I2C_Configuration.export
		.i2c_sdat        (trdb_d5m_camera_0_i2c_configuration_sdat), //                  .export
		.iexposure_adj   (trdb_d5m_camera_0_exposure_adjust_adj),    //   Exposure_Adjust.export
		.iexposure_dec_p (trdb_d5m_camera_0_exposure_adjust_dec_p),  //                  .export
		.iclk            (clk_clk),                                  //         iCLK_sink.clk
		.oRST_0          (trdb_d5m_camera_0_orst_0_reset),           //            oRST_0.reset
		.oRST_2          (trdb_d5m_camera_0_orst_2_reset),           //            oRST_2.reset
		.oRST_1          (trdb_d5m_camera_0_orst_1_reset),           //            oRST_1.reset
		.CCD_PIXCLK      (trdb_d5m_camera_0_ccd_pixclk_clk),         //        CCD_PIXCLK.clk
		.idata           (trdb_d5m_camera_0_idata_export),           //             idata.export
		.iend            (trdb_d5m_camera_0_iend_export),            //              iend.export
		.ifval           (trdb_d5m_camera_0_iflval_ifval),           //            iflval.export
		.ilval           (trdb_d5m_camera_0_iflval_ilval),           //                  .export
		.irst            (rst_controller_reset_out_reset),           //              irst.reset
		.istart          (trdb_d5m_camera_0_istart_export),          //            istart.export
		.izoom_mode_sw   (trdb_d5m_camera_0_zoom_mode_export),       //         zoom_mode.export
		.ored            (trdb_d5m_camera_0_rgb_ored),               //               rgb.export
		.ogreen          (trdb_d5m_camera_0_rgb_ogreen),             //                  .export
		.oblue           (trdb_d5m_camera_0_rgb_oblue),              //                  .export
		.odval           (trdb_d5m_camera_0_odval_export),           //             odval.export
		.oycont          (trdb_d5m_camera_0_oycont_export),          //            oycont.export
		.oframe          (trdb_d5m_camera_0_oframe_export)           //            oframe.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

endmodule
